module Decoder38(in, out);
input[2 : 0] in;
output[7 : 0] out;
assign out = 
	in == 0 ? 8'b00000001 : 
	in == 1 ? 8'b00000010 : 
	in == 2 ? 8'b00000100 : 
	in == 3 ? 8'b00001000 : 
	in == 4 ? 8'b00010000 : 
	in == 5 ? 8'b00100000 : 
	in == 6 ? 8'b01000000 : 
	in == 7 ? 8'b10000000 : 
	0;
endmodule

module Decode532(in, out);
input[4 : 0] in;
output[31 : 0] out;
assign out = 
	in == 0 ? 32'b00000000000000000000000000000001 : 
	in == 1 ? 32'b00000000000000000000000000000010 : 
	in == 2 ? 32'b00000000000000000000000000000100 : 
	in == 3 ? 32'b00000000000000000000000000001000 : 
	in == 4 ? 32'b00000000000000000000000000010000 : 
	in == 5 ? 32'b00000000000000000000000000100000 : 
	in == 6 ? 32'b00000000000000000000000001000000 : 
	in == 7 ? 32'b00000000000000000000000010000000 : 
	in == 8 ? 32'b00000000000000000000000100000000 : 
	in == 9 ? 32'b00000000000000000000001000000000 : 
	in == 10 ? 32'b00000000000000000000010000000000 : 
	in == 11 ? 32'b00000000000000000000100000000000 : 
	in == 12 ? 32'b00000000000000000001000000000000 : 
	in == 13 ? 32'b00000000000000000010000000000000 : 
	in == 14 ? 32'b00000000000000000100000000000000 : 
	in == 15 ? 32'b00000000000000001000000000000000 : 
	in == 16 ? 32'b00000000000000010000000000000000 : 
	in == 17 ? 32'b00000000000000100000000000000000 : 
	in == 18 ? 32'b00000000000001000000000000000000 : 
	in == 19 ? 32'b00000000000010000000000000000000 : 
	in == 20 ? 32'b00000000000100000000000000000000 : 
	in == 21 ? 32'b00000000001000000000000000000000 : 
	in == 22 ? 32'b00000000010000000000000000000000 : 
	in == 23 ? 32'b00000000100000000000000000000000 : 
	in == 24 ? 32'b00000001000000000000000000000000 : 
	in == 25 ? 32'b00000010000000000000000000000000 : 
	in == 26 ? 32'b00000100000000000000000000000000 : 
	in == 27 ? 32'b00001000000000000000000000000000 : 
	in == 28 ? 32'b00010000000000000000000000000000 : 
	in == 29 ? 32'b00100000000000000000000000000000 : 
	in == 30 ? 32'b01000000000000000000000000000000 : 
	in == 31 ? 32'b10000000000000000000000000000000 : 
0;
endmodule